1451624400,61832,
1454302800,64804,
1456808400,67816,
1459483200,71352,
1462075200,74690,
1464753600,77953,
1467345600,80832,1
1470024000,84063,2
1472702400,87398,3
1475294400,90619,4
1477972800,94001,5
1480568400,92745,
1483246800,95801,
1485925200,98785,
1488344400,102237,
1491019200,105977,
1493611200,109508,1
1496289600,104636,
1498881600,108017,
1501560000,111481,
1504238400,114802,
1506830400,117847,
1509508800,121412,1
1512104400,124960,2
1514782800,128414,3
1517461200,132457,4
1519880400,136051,5
1522555200,139820,6
1525147200,143609,7
1527825600,147383,8
1530417600,151403,9
1533096000,155355,10
1535774400,160660,11
1538366400,164469,12
1541044800,168440,13
1543640400,172797,14
1546318800,176355,15
1548997200,180653,16
1551416400,184829,17
1554091200,189569,18
1556683200,193991,19
1559361600,198698,20
1561953600,202758,21
1564632000,207139,22
1567310400,211522,23
1569902400,215907,24
1572580800,220080,25
1575176400,224194,26
1577854800,228405,27
1580533200,232761,28
1583038800,236650,29
1585713600,241107,30
1588305600,245775,31
1590984000,250628,32
1593576000,254765,33
1596254400,259175,34
1598932800,263389,35
1601524800,267518,36
1604203200,271635,37
1606798800,275613,38
1609477200,249683,
1612155600,253724,
1614574800,257382,
1617249600,263533,
1619841600,268668,
1622520000,273279,1

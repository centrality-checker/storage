1569902400,884722,
1572580800,888604,
1575176400,892738,
1577854800,896816,
1580533200,901201,
1583038800,905263,
1585713600,910135,1
1588305600,915009,2
1590984000,920185,3
1593576000,924939,4
1596254400,929887,5
1598932800,934775,6
1601524800,939761,7
1604203200,945235,8
1606798800,951454,9

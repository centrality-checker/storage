1328072400,4514,
1330578000,4672,
1333252800,4846,
1335844800,5041,
1338523200,5269,
1341115200,5505,
1343793600,5739,1
1346472000,6088,2
1349064000,6409,3
1351742400,6776,4
1354338000,7178,5
1357016400,7568,6
1359694800,8101,7
1362114000,8597,8
1364788800,9336,9
1367380800,10036,10
1370059200,10682,11
1372651200,11475,12
1375329600,12251,13
1378008000,12949,14
1380600000,13873,15
1383278400,14690,16
1385874000,15651,17
1388552400,16678,18
1391230800,17843,19
1393650000,18915,20
1396324800,20279,21
1398916800,21554,22
1401595200,22999,23
1404187200,24428,24
1406865600,25820,25
1409544000,27504,26
1412136000,29068,27
1414814400,30731,28
1417410000,32395,29
1420088400,33936,30
1422766800,35811,31
1425186000,37582,32
1427860800,39461,33
1430452800,41321,34
1433131200,43492,35
1435723200,45580,36
1438401600,48105,37
1441080000,50658,38
1443672000,53354,39
1446350400,56026,40
1448946000,58856,41
1451624400,61932,42
1454302800,64916,43
1456808400,67925,44
1459483200,71475,45
1462075200,74794,46
1464753600,78072,47
1467345600,80956,48
1470024000,84191,49
1472702400,87543,50
1475294400,90790,51
1477972800,94187,52
1480568400,92944,0
1483246800,96022,0
1485925200,99032,0
1488344400,102499,0
1491019200,106253,0
1493611200,109778,1
1496289600,104900,0
1498881600,108306,0
1501560000,111812,0
1504238400,115133,0
1506830400,118208,0
1509508800,121831,1
1512104400,125417,2
1514782800,128921,3
1517461200,132986,4
1519880400,136593,5
1522555200,140419,6
1525147200,144252,7
1527825600,148028,8
1530417600,152088,9
1533096000,156078,10
1535774400,161376,11
1538366400,165217,12
1541044800,169240,13
1543640400,173646,14
1546318800,177213,15
1548997200,181556,16
1551416400,185775,17
1554091200,190513,18
1556683200,195153,19
1559361600,199917,20
1561953600,204049,21
1564632000,208512,22
1567310400,212927,23
1569902400,217359,24
1572580800,221584,25
1575176400,225739,26
1577854800,229976,27
1580533200,234388,28
1583038800,238434,29
1585713600,243031,30
1588305600,247854,31
1590984000,252846,32
1593576000,257092,33
1596254400,261716,34
1598932800,266165,35
1601524800,270449,36
1604203200,275581,37
1606798800,281383,38
